library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_BRANCHING_PACKAGE.all;

--  THIS IS THE MAIN DRIVER FILE. 
	
ENTITY SEFA_MAIN IS
PORT (
		SEFA_IR_REGISTER_VALUE : IN STD_LOGIC_VECTOR(31 DOWNTO 0); 
		SEFA_clk : in std_logic; 
		SEFA_UPDATED_PC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_MAIN;


ARCHITECTURE arch OF SEFA_MAIN IS
	
	SIGNAL SEFA_OPCODE : STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL SEFA_RS_REGISTER_ADDRESS : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL SEFA_RT_REGISTER_ADDRESS : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL SEFA_IMMEDIATE16_VALUE : STD_LOGIC_VECTOR(15 DOWNTO 0); --BEQ BNE
	SIGNAL SEFA_IMMEDIATE26_VALUE : STD_LOGIC_VECTOR(25 DOWNTO 0); -- JUMP
	SIGNAL SEFA_RS_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_RT_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_CURRENT_PC_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_UPDATED_PC_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
BEGIN

	GET_IR_VALUES: SEFA_IR_REGISTER_DRIVER PORT MAP (
		SEFA_clk => SEFA_clk,
		SEFA_IR_REGISTER_VALUE => SEFA_IR_REGISTER_VALUE, 
		SEFA_OPCODE => SEFA_OPCODE,
		SEFA_RS_REGISTER_ADDRESS => SEFA_RS_REGISTER_ADDRESS, 
		SEFA_RT_REGISTER_ADDRESS => SEFA_RT_REGISTER_ADDRESS,
		SEFA_IMMEDIATE16_VALUE => SEFA_IMMEDIATE16_VALUE,
		SEFA_IMMEDIATE26_VALUE => SEFA_IMMEDIATE26_VALUE
		);
		
	GET_RS_RT_PC_VALUES: SEFA_REGISTER_MEMORY_FILE PORT MAP (
		SEFA_clk => SEFA_clk,
		SEFA_RS_REGISTER_ADDRESS => SEFA_RS_REGISTER_ADDRESS,
		SEFA_RT_REGISTER_ADDRESS => SEFA_RT_REGISTER_ADDRESS,
		SEFA_RS_VALUE => SEFA_RS_VALUE,
		SEFA_RT_VALUE => SEFA_RT_VALUE,
		SEFA_CURRENT_PC_VALUE => SEFA_CURRENT_PC_VALUE
		
	);
	
	
	
	NAL_CONTROLLER_AND_CONDITION: SEFA_COMPUTE_NAL_FROM_IR_VAL PORT MAP (
		SEFA_OPCODE => SEFA_OPCODE,
		SEFA_RS_VALUE => SEFA_RS_VALUE,
		SEFA_RT_VALUE => SEFA_RT_VALUE, 
		SEFA_PC_VALUE => SEFA_CURRENT_PC_VALUE,
		SEFA_IMM16_VAL => SEFA_IMMEDIATE16_VALUE,
		SEFA_IMM26_VAL => SEFA_IMMEDIATE26_VALUE,
		SEFA_UPDATED_PC => SEFA_UPDATED_PC_VALUE
		
	);

	
	SEFA_UPDATED_PC <= SEFA_UPDATED_PC_VALUE; 
	
	
	


END arch; 

