library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_BRANCHING_PACKAGE.all;


ENTITY SEFA_BRANCHING_SIGNED_EXTENDED IS
PORT(
		
		SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		SEFA_SIGNED_16_to_32_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_SIGNED_26_to_32_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_SIGNED_32_EXTENDED_IMM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_BRANCHING_SIGNED_EXTENDED;

ARCHITECTURE arch OF SEFA_BRANCHING_SIGNED_EXTENDED IS
	
BEGIN


	SEFA_SIGNED_32_EXTENDED_IMM <= SEFA_SIGNED_26_to_32_EXTENDED_IMM WHEN SEFA_OPCODE = "111111"
							ELSE SEFA_SIGNED_16_to_32_EXTENDED_IMM;

END arch;
