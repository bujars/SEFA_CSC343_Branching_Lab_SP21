library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_BRANCHING_PACKAGE.all;



ENTITY SEFA_COMPUTE_NAL_FROM_IR_VAL IS 
PORT(
	
	
	
	 RS_VALUE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	 RT_VALUE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	 PC_VALUE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	 IMM16_VAL : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	SEFA_PC_NEW : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)  
);
END SEFA_COMPUTE_NAL_FROM_IR_VAL;


ARCHITECTURE arch OF SEFA_COMPUTE_NAL_FROM_IR_VAL IS

-- comparator value
	SIGNAL PC_COND : STD_LOGIC;

-- TO GET RESULT SO WE CAN STORE INTO RAM. 
	SIGNAL PC_UPDATED : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
	
	
	-- AFTER GETTING RS AND RT, COMPARE THEIR VALUES TO SET CONDITION
	COMPUTE_RS_RT_COMPARE : SEFA_Comparator_N PORT MAP (
		SEFA_IN0 => RS_VALUE, 
	
	SEFA_IN1 => RT_VALUE,
		SEFA_OUT => PC_COND
	
	);
	
	-- USING CONDITION AND PC, UPDATE THE NEW PC.
	COMPUTE_NAL : SEFA_NAL PORT MAP (
		SEFA_PC_COND => PC_COND, 
		SEFA_PC_OLD => PC_VALUE,
		SEFA_IMM16 => IMM16_VAL,
		SEFA_PC_NEW_OUT => SEFA_PC_NEW
	);

END arch; 