library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_BRANCHING_PACKAGE.all;



ENTITY SEFA_COMPUTE_NAL_FROM_IR_VAL IS 
PORT(
	 SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	 SEFA_RS_VALUE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	 SEFA_RT_VALUE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	 SEFA_PC_VALUE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	 SEFA_IMM16_VAL : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	 SEFA_IMM26_VAL : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
	 SEFA_UPDATED_PC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)  
	 
);
END SEFA_COMPUTE_NAL_FROM_IR_VAL;


ARCHITECTURE arch OF SEFA_COMPUTE_NAL_FROM_IR_VAL IS

-- comparator value
	SIGNAL SEFA_PC_COND : STD_LOGIC;

-- TO GET RESULT SO WE CAN STORE INTO RAM. 
	SIGNAL PC_UPDATED : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
	
	
	-- AFTER GETTING RS AND RT, COMPARE THEIR VALUES TO SET CONDITION
	COMPUTE_RS_RT_COMPARE : SEFA_Comparator_N PORT MAP (
		SEFA_IN0 => SEFA_RS_VALUE, 
	
	SEFA_IN1 => SEFA_RT_VALUE,
		SEFA_OUT => SEFA_PC_COND
	
	);
	
	
	-- ^ THIS WONT MATTER FOR JUMP!
	
	
	-- USING CONDITION AND PC, UPDATE THE NEW PC.
	COMPUTE_NAL : SEFA_NAL PORT MAP (
		SEFA_OPCODE => SEFA_OPCODE, 
		SEFA_PC_COND => SEFA_PC_COND, 
		SEFA_PC_OLD => SEFA_PC_VALUE,
		SEFA_IMM16 => SEFA_IMM16_VAL,
		SEFA_IMM26 => SEFA_IMM26_VAL,
		SEFA_UPDATED_PC => SEFA_UPDATED_PC
	);

END arch; 