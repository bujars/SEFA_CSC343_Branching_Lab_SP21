library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_BRANCHING_PACKAGE.all;

-- THE PURPOSE OF THIS COMPONENT IS TO SET THE FIELDS
-- OF DATA
-- THAT IS OPCODE | RS | RT | IMM16
-- we also might be able to avoid this file and do ir directly in IR_register
-- but im using ir register just for the sake of storing (read/write) data

ENTITY SEFA_IR_REGISTER_DRIVER IS
PORT (
	SEFA_clk: in std_logic;
	SEFA_IR_REGISTER_VALUE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	 SEFA_OPCODE : OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
	 SEFA_RS_REGISTER_ADDRESS : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
	 SEFA_RT_REGISTER_ADDRESS : OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
	 SEFA_IMMEDIATE16_VALUE : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	 SEFA_IMMEDIATE26_VALUE : OUT STD_LOGIC_VECTOR(25 DOWNTO 0)
);
END SEFA_IR_REGISTER_DRIVER;

ARCHITECTURE arch OF SEFA_IR_REGISTER_DRIVER IS
	SIGNAL SEFA_IR_REGISTER_VALUE_OUTPUT: STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN


	SET_AND_GET_IR_VALUE_IN_REGISTER : SEFA_IR_REGISTER port map (
		SEFA_clk => SEFA_clk, 
		SEFA_wren => '1',
		SEFA_rden => '1', 
		SEFA_chen => '1', 
		SEFA_data => SEFA_IR_REGISTER_VALUE, 
		SEFA_IR=> SEFA_IR_REGISTER_VALUE_OUTPUT
	);
	

	SEFA_OPCODE <= SEFA_IR_REGISTER_VALUE_OUTPUT(31 DOWNTO 26);
	SEFA_RS_REGISTER_ADDRESS <= SEFA_IR_REGISTER_VALUE_OUTPUT(25 DOWNTO 21);
	SEFA_RT_REGISTER_ADDRESS <= SEFA_IR_REGISTER_VALUE_OUTPUT(20 DOWNTO 16);
	SEFA_IMMEDIATE16_VALUE <= SEFA_IR_REGISTER_VALUE_OUTPUT(15 DOWNTO 0);
	
	
	
	-- NOTE. WHEN JUMP IS EXECUTING, THE RESUT OF THE VALUES WILL HAVE "JUNK" 
	-- WHEN EXECUTING RS RT IMM16, WELL THOSE ARE SIMPLY STORED IN IMM26 (BUT WE WONT USE IT)
	SEFA_IMMEDIATE26_VALUE <= SEFA_IR_REGISTER_VALUE_OUTPUT(25 DOWNTO 0);

	


END arch;

