library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_BRANCHING_PACKAGE.all;


-- NOTE THIS FILE ESSENTIALLY REPLACES THE MUX
-- THIS IS BECAUSE WE WANT TO SIMPLFY THE LOGIC OF COMPUTING TEH ADDRESSES
-- IE COMPUTE BASED ON CONDITION, NOT COMPUTE AND THEN SELECT THE GIVEN RESULT. 
-- THIS IS SIMILAR TO THE ORIGINAL ERROR MADE IN LAB1 BUT THEN YOU CORRECTED IT. 
-- IT WILL REQUIRE A IF-ELSE (WITH PROCESS)

-- had to go select result. Compute on condition does not seem to be working for me. Maybe im misunderstanding what can go in if...


ENTITY SEFA_NAL IS
PORT(
		SEFA_PC_COND : IN STD_LOGIC;
		SEFA_PC_OLD : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_IMM16 : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- NOTE THIS IS 16 BITS AND WE NEED TO SIGN EXTEND! 
		SEFA_PC_NEW_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_NAL;

ARCHITECTURE arch OF SEFA_NAL IS

	SIGNAL SIGNED_EXTENDED_IMM : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_PLUS_4 : STD_LOGIC_VECTOR(31 DOWNTO 0); -- NOTE THIS IS NEEDED FOR EITHER MODULE, SO ITS COMPUTED IN THE BEGINNING
	SIGNAL PC_PLUS_IMM_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	
BEGIN
	
	PC_4: SEFA_PC_PLUS_4 PORT MAP (
						SEFA_PC_OLD => SEFA_PC_OLD,
						SEFA_PC_NEW => PC_PLUS_4
	);
	
	A: SEFA_SIGN_EXTEND_IMM_16_TO_32 PORT MAP ( SEFA_IMM16 => SEFA_IMM16, SEFA_IMM32 => SIGNED_EXTENDED_IMM);
	B: SEFA_PC_PLUS_IMMEDIATE_PLUS_4 PORT MAP ( SEFA_PC_PLUS_4 => PC_PLUS_4, SEFA_SIGN_EXTENDED_IMM => SIGNED_EXTENDED_IMM, SEFA_PC_NEW => PC_PLUS_IMM_4 );	
	
--	
--	PROCESS (SEFA_PC_COND)
--	BEGIN
--	
--		-- HANDLE JUMPING VIA IMMEDIATE
--		IF (SEFA_PC_COND = '1') THEN
--				SEFA_PC_NEW_OUT <= PC_PLUS_IMM_4;
--		ELSE -- CONTINUE TO NEXT ADDRESS (+4)
--			SEFA_PC_NEW_OUT <= PC_PLUS_4;
--		END IF;
--	
--	END PROCESS;
	C: SEFA_Branching_MUX PORT MAP ( SEFA_PC_Plus_4 =>  PC_PLUS_4, SEFA_PC_IMM16_Plus_4 => PC_PLUS_IMM_4, SEFA_PC_SELECTOR => SEFA_PC_COND, SEFA_PC_NEW => SEFA_PC_NEW_OUT);

END arch;