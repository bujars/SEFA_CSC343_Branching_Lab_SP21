library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_BRANCHING_PACKAGE.all;


-- NOTE THIS FILE ESSENTIALLY REPLACES THE MUX
-- THIS IS BECAUSE WE WANT TO SIMPLFY THE LOGIC OF COMPUTING TEH ADDRESSES
-- IE COMPUTE BASED ON CONDITION, NOT COMPUTE AND THEN SELECT THE GIVEN RESULT. 
-- THIS IS SIMILAR TO THE ORIGINAL ERROR MADE IN LAB1 BUT THEN YOU CORRECTED IT. 
-- IT WILL REQUIRE A IF-ELSE (WITH PROCESS)

ENTITY SEFA_NAL IS
PORT(
		SEFA_PC_COND : IN STD_LOGIC;
		SEFA_PC_OLD : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_IMM16 : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- NOTE THIS IS 16 BITS AND WE NEED TO SIGN EXTEND! 
		SEFA_PC_NEW : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
);
END SEFA_NAL;

ARCHITECTURE arch OF SEFA_NAL IS

SIGNAL SEFA_SIGNED_EXTENDED_IMM : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL SEFA_PC_PLUS_4 : STD_LOGIC_VECTOR(31 DOWNTO 0); -- NOTE THIS IS NEEDED FOR EITHER MODULE, SO ITS COMPUTED IN THE BEGINNING

BEGIN
	
	SEFA_PC_PLUS_4: SEFA_PC_PLUS_4 PORT MAP (
						SEFA_PC_OLD => SEFA_PC_OLD,
						SEFA_PC_NEW => SEFA_PC_PLUS_4
	);

	PROCESS(SEFA_PC_COND, SEFA_PC_OLD, SEFA_IMM16)
	BEGIN
	
		-- HANDLE JUMPING VIA IMMEDIATE
		IF (SEFA_PC_COND = 1) THEN
			SIGNED_EXTENDED: SEFA_SIGN_EXTEND_IMM_16_TO_32 PORT MAP (
						SEFA_IMM16 => SEFA_IMM16,
						SEFA_IMM32 => SEFA_SIGNED_EXTENDED_IMM
			);
			PC_PLUS_4_PLUS_IMMEDIATE: SEFA_PC_PLUS_IMMEDIATE_PLUS_4 PORT MAP (
						SEFA_PC_PLUS_4 => SEFA_PC_PLUS_4,
						SEFA_SIGN_EXTENDED_IMM => SEFA_SIGNED_EXTENDED_IMM,
						SEFA_PC_NEW => SEFA_PC_NEW
			);	
		ELSE -- CONTINUE TO NEXT ADDRESS (+4)
			SEFA_PC_NEW <= SEFA_PC_PLUS_4;
		
		END IF;
	
	END PROCESS;

END arch;