library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_BRANCHING_PACKAGE.all;

-- SEFA_REGISTER_MEMORY_FILE

ENTITY SEFA_REGISTER_MEMORY_FILE IS 
PORT  
(
		SEFA_clk : IN STD_LOGIC; 
		SEFA_RS_REGISTER_ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		SEFA_RT_REGISTER_ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		SEFA_RS_VALUE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_RT_VALUE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_CURRENT_PC_VALUE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		
	);
END SEFA_REGISTER_MEMORY_FILE;

ARCHITECTURE arch OF SEFA_REGISTER_MEMORY_FILE IS

	SIGNAL SEFA_RS_MEMORY_OUTPUT_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_RT_MEMORY_OUTPUT_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_CURRENT_PC_MEMORY_OUTPUT_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
--	SIGNAL SEFA_RS_REGISTER_OUTPUT_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
--	SIGNAL SEFA_RT_REGISTER_OUTPUT_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
--	SIGNAL SEFA_CURRENT_PC_REGISTER_OUTPUT_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
	GET_PC_VALUE_FROM_MEMORY: SEFA_INSTRUCTION_MEMORY PORT MAP (
		address => "00000", -- THE PC IS default address HERE! MUST BE CONSISTENT ON ALL FILES THAT PULL IT OR NEED THE ADDRESS. 
		clock => SEFA_clk,
		data => "00000000000000000000000000000000", -- arbitrary because we are reading
		wren => '0',
		q => SEFA_CURRENT_PC_MEMORY_OUTPUT_VALUE
		
	);
	
	GET_RS_VALUE_FROM_MEMORY: SEFA_INSTRUCTION_MEMORY PORT MAP (
		address => SEFA_RS_REGISTER_ADDRESS,
		clock => SEFA_clk,
		data => "00000000000000000000000000000000", -- NOTE THIS IS ANY ARBITRARY DATA BECAUSE WE AREN'T WRITING TO IT. ONLY READING RS!
		wren => '0',
		q => SEFA_RS_MEMORY_OUTPUT_VALUE
	);
	
	GET_RT_VALUE_MEMORY: SEFA_INSTRUCTION_MEMORY PORT MAP (
		address => SEFA_RT_REGISTER_ADDRESS,
		clock => SEFA_clk,
		data => "00000000000000000000000000000000", -- NOTE THIS IS ANY ARBITRARY DATA BECAUSE WE AREN'T WRITING TO IT. ONLY READING RT!
		wren => '0',
		q => SEFA_RT_MEMORY_OUTPUT_VALUE
	);

	SET_AND_GET_PC_VALUE_IN_REGISTER : SEFA_PC_REGISTER port map (
		SEFA_clk => SEFA_clk, 
		SEFA_wren => '1',
		SEFA_rden => '1', 
		SEFA_chen => '1', 
		SEFA_data => SEFA_CURRENT_PC_MEMORY_OUTPUT_VALUE, 
		SEFA_PC=> SEFA_CURRENT_PC_VALUE
	);
	
	SET_AND_GET_RS_VALUE_IN_REGISTER : SEFA_RS_REGISTER port map (
		SEFA_clk => SEFA_clk, 
		SEFA_wren => '1',
		SEFA_rden => '1', 
		SEFA_chen => '1', 
		SEFA_data => SEFA_RS_MEMORY_OUTPUT_VALUE, 
		SEFA_RS=> SEFA_RS_VALUE
	);
	
	SET_AND_GET_RT_VALUE_IN_REGISTER : SEFA_RT_REGISTER port map (
		SEFA_clk => SEFA_clk, 
		SEFA_wren => '1',
		SEFA_rden => '1', 
		SEFA_chen => '1', 
		SEFA_data => SEFA_RT_MEMORY_OUTPUT_VALUE, 
		SEFA_RT=> SEFA_RT_VALUE
	);





END arch;